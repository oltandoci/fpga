-- BRIEF    : Project configuration
-- DATE     : March 23th, 2015
-- AUTHOR   : O.D

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE proj_config IS

    CONSTANT C_MEM_POWER_2_DEPTH    : POSITIVE := 8; --Number of FFT samples = 2^C_MEM_POWER_2_DEPTH i.e. 256 here
    CONSTANT C_MEM_DATA_LENGTH      : POSITIVE := 16;
    CONSTANT C_CRC_POLYNOMIAL32     : STD_LOGIC_VECTOR(31 DOWNTO 0) := X"04C11DB7";
    
    TYPE t_sin_cos_table IS ARRAY (0 TO ((2**C_MEM_POWER_2_DEPTH) - 1)) OF STD_LOGIC_VECTOR(C_MEM_DATA_LENGTH - 1 DOWNTO 0);
    TYPE t_crc_table IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR(15 DOWNTO 0);

END PACKAGE proj_config;
